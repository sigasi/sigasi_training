library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity dummy is -- TODO: delete this file
	port (
		clk : in std_logic;
		rst : in std_logic
	);
end entity dummy;
