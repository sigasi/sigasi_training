library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity dummy is
	port (
		clk : in std_logic;
		rst : in std_logic
	);
end entity dummy;

architecture RTL of dummy is
	
begin
	
end architecture RTL;

