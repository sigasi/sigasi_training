library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity duplicate is
	port (
		clk : in std_logic;
		rst : in std_logic
	);
end entity duplicate;
